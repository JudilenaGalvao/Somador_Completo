library verilog;
use verilog.vl_types.all;
entity SomadorCompleto_vlg_vec_tst is
end SomadorCompleto_vlg_vec_tst;
